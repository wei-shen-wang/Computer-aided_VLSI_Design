module sq(
    input [7:0] sq_in, //s1.6
    input sq_en,
    output reg [7:0] sq_out //0.8
);
    

    always@(*) begin

        if (sq_en) begin
        case(sq_in)

        default : sq_out = 8'b11111111;

        8'b00000000 : sq_out = 8'b00000000;
        8'b00000001 : sq_out = 8'b00000000;
        8'b00000010 : sq_out = 8'b00000000;
        8'b00000011 : sq_out = 8'b00000001;
        8'b00000100 : sq_out = 8'b00000001;
        8'b00000101 : sq_out = 8'b00000010;
        8'b00000110 : sq_out = 8'b00000010;
        8'b00000111 : sq_out = 8'b00000011;
        8'b00001000 : sq_out = 8'b00000100;
        8'b00001001 : sq_out = 8'b00000101;
        8'b00001010 : sq_out = 8'b00000110;
        8'b00001011 : sq_out = 8'b00001000;
        8'b00001100 : sq_out = 8'b00001001;
        8'b00001101 : sq_out = 8'b00001011;
        8'b00001110 : sq_out = 8'b00001100;
        8'b00001111 : sq_out = 8'b00001110;
        8'b00010000 : sq_out = 8'b00010000;
        8'b00010001 : sq_out = 8'b00010010;
        8'b00010010 : sq_out = 8'b00010100;
        8'b00010011 : sq_out = 8'b00010111;
        8'b00010100 : sq_out = 8'b00011001;
        8'b00010101 : sq_out = 8'b00011100;
        8'b00010110 : sq_out = 8'b00011110;
        8'b00010111 : sq_out = 8'b00100001;
        8'b00011000 : sq_out = 8'b00100100;
        8'b00011001 : sq_out = 8'b00100111;
        8'b00011010 : sq_out = 8'b00101010;
        8'b00011011 : sq_out = 8'b00101110;
        8'b00011100 : sq_out = 8'b00110001;
        8'b00011101 : sq_out = 8'b00110101;
        8'b00011110 : sq_out = 8'b00111000;
        8'b00011111 : sq_out = 8'b00111100;
        8'b00100000 : sq_out = 8'b01000000;
        8'b00100001 : sq_out = 8'b01000100;
        8'b00100010 : sq_out = 8'b01001000;
        8'b00100011 : sq_out = 8'b01001101;
        8'b00100100 : sq_out = 8'b01010001;
        8'b00100101 : sq_out = 8'b01010110;
        8'b00100110 : sq_out = 8'b01011010;
        8'b00100111 : sq_out = 8'b01011111;
        8'b00101000 : sq_out = 8'b01100100;
        8'b00101001 : sq_out = 8'b01101001;
        8'b00101010 : sq_out = 8'b01101110;
        8'b00101011 : sq_out = 8'b01110100;
        8'b00101100 : sq_out = 8'b01111001;
        8'b00101101 : sq_out = 8'b01111111;
        8'b00101110 : sq_out = 8'b10000100;
        8'b00101111 : sq_out = 8'b10001010;
        8'b00110000 : sq_out = 8'b10010000;
        8'b00110001 : sq_out = 8'b10010110;
        8'b00110010 : sq_out = 8'b10011100;
        8'b00110011 : sq_out = 8'b10100011;
        8'b00110100 : sq_out = 8'b10101001;
        8'b00110101 : sq_out = 8'b10110000;
        8'b00110110 : sq_out = 8'b10110110;
        8'b00110111 : sq_out = 8'b10111101;
        8'b00111000 : sq_out = 8'b11000100;
        8'b00111001 : sq_out = 8'b11001011;
        8'b00111010 : sq_out = 8'b11010010;
        8'b00111011 : sq_out = 8'b11011010;
        8'b00111100 : sq_out = 8'b11100001;
        8'b00111101 : sq_out = 8'b11101001;
        8'b00111110 : sq_out = 8'b11110000;
        8'b00111111 : sq_out = 8'b11111000;

        8'b11000001 : sq_out = 8'b11111000;
        8'b11000010 : sq_out = 8'b11110000;
        8'b11000011 : sq_out = 8'b11101001;
        8'b11000100 : sq_out = 8'b11100001;
        8'b11000101 : sq_out = 8'b11011010;
        8'b11000110 : sq_out = 8'b11010010;
        8'b11000111 : sq_out = 8'b11001011;
        8'b11001000 : sq_out = 8'b11000100;
        8'b11001001 : sq_out = 8'b10111101;
        8'b11001010 : sq_out = 8'b10110110;
        8'b11001011 : sq_out = 8'b10110000;
        8'b11001100 : sq_out = 8'b10101001;
        8'b11001101 : sq_out = 8'b10100011;
        8'b11001110 : sq_out = 8'b10011100;
        8'b11001111 : sq_out = 8'b10010110;
        8'b11010000 : sq_out = 8'b10010000;
        8'b11010001 : sq_out = 8'b10001010;
        8'b11010010 : sq_out = 8'b10000100;
        8'b11010011 : sq_out = 8'b01111111;
        8'b11010100 : sq_out = 8'b01111001;
        8'b11010101 : sq_out = 8'b01110100;
        8'b11010110 : sq_out = 8'b01101110;
        8'b11010111 : sq_out = 8'b01101001;
        8'b11011000 : sq_out = 8'b01100100;
        8'b11011001 : sq_out = 8'b01011111;
        8'b11011010 : sq_out = 8'b01011010;
        8'b11011011 : sq_out = 8'b01010110;
        8'b11011100 : sq_out = 8'b01010001;
        8'b11011101 : sq_out = 8'b01001101;
        8'b11011110 : sq_out = 8'b01001000;
        8'b11011111 : sq_out = 8'b01000100;
        8'b11100000 : sq_out = 8'b01000000;
        8'b11100001 : sq_out = 8'b00111100;
        8'b11100010 : sq_out = 8'b00111000;
        8'b11100011 : sq_out = 8'b00110101;
        8'b11100100 : sq_out = 8'b00110001;
        8'b11100101 : sq_out = 8'b00101110;
        8'b11100110 : sq_out = 8'b00101010;
        8'b11100111 : sq_out = 8'b00100111;
        8'b11101000 : sq_out = 8'b00100100;
        8'b11101001 : sq_out = 8'b00100001;
        8'b11101010 : sq_out = 8'b00011110;
        8'b11101011 : sq_out = 8'b00011100;
        8'b11101100 : sq_out = 8'b00011001;
        8'b11101101 : sq_out = 8'b00010111;
        8'b11101110 : sq_out = 8'b00010100;
        8'b11101111 : sq_out = 8'b00010010;
        8'b11110000 : sq_out = 8'b00010000;
        8'b11110001 : sq_out = 8'b00001110;
        8'b11110010 : sq_out = 8'b00001100;
        8'b11110011 : sq_out = 8'b00001011;
        8'b11110100 : sq_out = 8'b00001001;
        8'b11110101 : sq_out = 8'b00001000;
        8'b11110110 : sq_out = 8'b00000110;
        8'b11110111 : sq_out = 8'b00000101;
        8'b11111000 : sq_out = 8'b00000100;
        8'b11111001 : sq_out = 8'b00000011;
        8'b11111010 : sq_out = 8'b00000010;
        8'b11111011 : sq_out = 8'b00000010;
        8'b11111100 : sq_out = 8'b00000001;
        8'b11111101 : sq_out = 8'b00000001;
        8'b11111110 : sq_out = 8'b00000000;
        8'b11111111 : sq_out = 8'b00000000;

        endcase
        end
        else sq_out = 0;

    end
endmodule