module sqrt(
    input [10:0] sqrt_in, //3.8
    output reg [19:0] sqrt_out //S3.16
);
    

    always@(*) begin
        casez(sqrt_in)

            default : sqrt_out = 20'b00000001000000000000;

            // 13'b1zzzzzzzzzzzz : sqrt_out = 20'b01000000000000000000;
            
            // 13'b01zzzzzzzzzzz : sqrt_out = 20'b00101101010000010011; 
            
            11'b10zzzzzzzzz : sqrt_out = 20'b00100000000000000000;
            11'b11zzzzzzzzz : sqrt_out = 20'b00100111001100010001;

            11'b010000000zz : sqrt_out = 20'b00010110101000001001;
            11'b010000001zz : sqrt_out = 20'b00010110101101110011;
            11'b010000010zz : sqrt_out = 20'b00010110110011011011;
            11'b010000011zz : sqrt_out = 20'b00010110111001000001;
            11'b010000100zz : sqrt_out = 20'b00010110111110100110;
            11'b010000101zz : sqrt_out = 20'b00010111000100001010;
            11'b010000110zz : sqrt_out = 20'b00010111001001101101;
            11'b010000111zz : sqrt_out = 20'b00010111001111001110;
            11'b010001000zz : sqrt_out = 20'b00010111010100101110;
            11'b010001001zz : sqrt_out = 20'b00010111011010001100;
            11'b010001010zz : sqrt_out = 20'b00010111011111101010;
            11'b010001011zz : sqrt_out = 20'b00010111100101000110;
            11'b010001100zz : sqrt_out = 20'b00010111101010100001;
            11'b010001101zz : sqrt_out = 20'b00010111101111111010;
            11'b010001110zz : sqrt_out = 20'b00010111110101010010;
            11'b010001111zz : sqrt_out = 20'b00010111111010101010;
            11'b010010000zz : sqrt_out = 20'b00011000000000000000;
            11'b010010001zz : sqrt_out = 20'b00011000000101010100;
            11'b010010010zz : sqrt_out = 20'b00011000001010101000;
            11'b010010011zz : sqrt_out = 20'b00011000001111111010;
            11'b010010100zz : sqrt_out = 20'b00011000010101001011;
            11'b010010101zz : sqrt_out = 20'b00011000011010011100;
            11'b010010110zz : sqrt_out = 20'b00011000011111101011;
            11'b010010111zz : sqrt_out = 20'b00011000100100111000;
            11'b010011000zz : sqrt_out = 20'b00011000101010000101;
            11'b010011001zz : sqrt_out = 20'b00011000101111010001;
            11'b010011010zz : sqrt_out = 20'b00011000110100011100;
            11'b010011011zz : sqrt_out = 20'b00011000111001100101;
            11'b010011100zz : sqrt_out = 20'b00011000111110101110;
            11'b010011101zz : sqrt_out = 20'b00011001000011110101;
            11'b010011110zz : sqrt_out = 20'b00011001001000111011;
            11'b010011111zz : sqrt_out = 20'b00011001001110000001;
            11'b010100000zz : sqrt_out = 20'b00011001010011000101;
            11'b010100001zz : sqrt_out = 20'b00011001011000001000;
            11'b010100010zz : sqrt_out = 20'b00011001011101001011;
            11'b010100011zz : sqrt_out = 20'b00011001100010001100;
            11'b010100100zz : sqrt_out = 20'b00011001100111001100;
            11'b010100101zz : sqrt_out = 20'b00011001101100001100;
            11'b010100110zz : sqrt_out = 20'b00011001110001001010;
            11'b010100111zz : sqrt_out = 20'b00011001110110000111;
            11'b010101000zz : sqrt_out = 20'b00011001111011000100;
            11'b010101001zz : sqrt_out = 20'b00011010000000000000;
            11'b010101010zz : sqrt_out = 20'b00011010000100111010;
            11'b010101011zz : sqrt_out = 20'b00011010001001110100;
            11'b010101100zz : sqrt_out = 20'b00011010001110101101;
            11'b010101101zz : sqrt_out = 20'b00011010010011100100;
            11'b010101110zz : sqrt_out = 20'b00011010011000011011;
            11'b010101111zz : sqrt_out = 20'b00011010011101010001;
            11'b010110000zz : sqrt_out = 20'b00011010100010000111;
            11'b010110001zz : sqrt_out = 20'b00011010100110111011;
            11'b010110010zz : sqrt_out = 20'b00011010101011101110;
            11'b010110011zz : sqrt_out = 20'b00011010110000100001;
            11'b010110100zz : sqrt_out = 20'b00011010110101010011;
            11'b010110101zz : sqrt_out = 20'b00011010111010000100;
            11'b010110110zz : sqrt_out = 20'b00011010111110110100;
            11'b010110111zz : sqrt_out = 20'b00011011000011100011;
            11'b010111000zz : sqrt_out = 20'b00011011001000010001;
            11'b010111001zz : sqrt_out = 20'b00011011001100111111;
            11'b010111010zz : sqrt_out = 20'b00011011010001101011;
            11'b010111011zz : sqrt_out = 20'b00011011010110010111;
            11'b010111100zz : sqrt_out = 20'b00011011011011000011;
            11'b010111101zz : sqrt_out = 20'b00011011011111101101;
            11'b010111110zz : sqrt_out = 20'b00011011100100010110;
            11'b010111111zz : sqrt_out = 20'b00011011101000111111;
            11'b011000000zz : sqrt_out = 20'b00011011101101100111;
            11'b011000001zz : sqrt_out = 20'b00011011110010001110;
            11'b011000010zz : sqrt_out = 20'b00011011110110110101;
            11'b011000011zz : sqrt_out = 20'b00011011111011011011;
            11'b011000100zz : sqrt_out = 20'b00011100000000000000;
            11'b011000101zz : sqrt_out = 20'b00011100000100100100;
            11'b011000110zz : sqrt_out = 20'b00011100001001000111;
            11'b011000111zz : sqrt_out = 20'b00011100001101101010;
            11'b011001000zz : sqrt_out = 20'b00011100010010001100;
            11'b011001001zz : sqrt_out = 20'b00011100010110101101;
            11'b011001010zz : sqrt_out = 20'b00011100011011001110;
            11'b011001011zz : sqrt_out = 20'b00011100011111101110;
            11'b011001100zz : sqrt_out = 20'b00011100100100001101;
            11'b011001101zz : sqrt_out = 20'b00011100101000101011;
            11'b011001110zz : sqrt_out = 20'b00011100101101001001;
            11'b011001111zz : sqrt_out = 20'b00011100110001100110;
            11'b011010000zz : sqrt_out = 20'b00011100110110000010;
            11'b011010001zz : sqrt_out = 20'b00011100111010011110;
            11'b011010010zz : sqrt_out = 20'b00011100111110111001;
            11'b011010011zz : sqrt_out = 20'b00011101000011010011;
            11'b011010100zz : sqrt_out = 20'b00011101000111101101;
            11'b011010101zz : sqrt_out = 20'b00011101001100000110;
            11'b011010110zz : sqrt_out = 20'b00011101010000011110;
            11'b011010111zz : sqrt_out = 20'b00011101010100110110;
            11'b011011000zz : sqrt_out = 20'b00011101011001001101;
            11'b011011001zz : sqrt_out = 20'b00011101011101100011;
            11'b011011010zz : sqrt_out = 20'b00011101100001111001;
            11'b011011011zz : sqrt_out = 20'b00011101100110001110;
            11'b011011100zz : sqrt_out = 20'b00011101101010100010;
            11'b011011101zz : sqrt_out = 20'b00011101101110110110;
            11'b011011110zz : sqrt_out = 20'b00011101110011001010;
            11'b011011111zz : sqrt_out = 20'b00011101110111011100;
            11'b011100000zz : sqrt_out = 20'b00011101111011101110;
            11'b011100001zz : sqrt_out = 20'b00011110000000000000;
            11'b011100010zz : sqrt_out = 20'b00011110000100010000;
            11'b011100011zz : sqrt_out = 20'b00011110001000100000;
            11'b011100100zz : sqrt_out = 20'b00011110001100110000;
            11'b011100101zz : sqrt_out = 20'b00011110010000111111;
            11'b011100110zz : sqrt_out = 20'b00011110010101001101;
            11'b011100111zz : sqrt_out = 20'b00011110011001011011;
            11'b011101000zz : sqrt_out = 20'b00011110011101101000;
            11'b011101001zz : sqrt_out = 20'b00011110100001110101;
            11'b011101010zz : sqrt_out = 20'b00011110100110000001;
            11'b011101011zz : sqrt_out = 20'b00011110101010001100;
            11'b011101100zz : sqrt_out = 20'b00011110101110010111;
            11'b011101101zz : sqrt_out = 20'b00011110110010100010;
            11'b011101110zz : sqrt_out = 20'b00011110110110101100;
            11'b011101111zz : sqrt_out = 20'b00011110111010110101;
            11'b011110000zz : sqrt_out = 20'b00011110111110111101;
            11'b011110001zz : sqrt_out = 20'b00011111000011000110;
            11'b011110010zz : sqrt_out = 20'b00011111000111001101;
            11'b011110011zz : sqrt_out = 20'b00011111001011010100;
            11'b011110100zz : sqrt_out = 20'b00011111001111011011;
            11'b011110101zz : sqrt_out = 20'b00011111010011100001;
            11'b011110110zz : sqrt_out = 20'b00011111010111100110;
            11'b011110111zz : sqrt_out = 20'b00011111011011101011;
            11'b011111000zz : sqrt_out = 20'b00011111011111101111;
            11'b011111001zz : sqrt_out = 20'b00011111100011110011;
            11'b011111010zz : sqrt_out = 20'b00011111100111110110;
            11'b011111011zz : sqrt_out = 20'b00011111101011111001;
            11'b011111100zz : sqrt_out = 20'b00011111101111111011;
            11'b011111101zz : sqrt_out = 20'b00011111110011111101;
            11'b011111110zz : sqrt_out = 20'b00011111110111111110;
            11'b011111111zz : sqrt_out = 20'b00011111111011111111;

            11'b00100000000 : sqrt_out = 20'b00010000000000000000;
            11'b00100000001 : sqrt_out = 20'b00010000000001111111;
            11'b00100000010 : sqrt_out = 20'b00010000000011111111;
            11'b00100000011 : sqrt_out = 20'b00010000000101111110;
            11'b00100000100 : sqrt_out = 20'b00010000000111111110;
            11'b00100000101 : sqrt_out = 20'b00010000001001111100;
            11'b00100000110 : sqrt_out = 20'b00010000001011111011;
            11'b00100000111 : sqrt_out = 20'b00010000001101111001;
            11'b00100001000 : sqrt_out = 20'b00010000001111111000;
            11'b00100001001 : sqrt_out = 20'b00010000010001110110;
            11'b00100001010 : sqrt_out = 20'b00010000010011110011;
            11'b00100001011 : sqrt_out = 20'b00010000010101110001;
            11'b00100001100 : sqrt_out = 20'b00010000010111101110;
            11'b00100001101 : sqrt_out = 20'b00010000011001101011;
            11'b00100001110 : sqrt_out = 20'b00010000011011101000;
            11'b00100001111 : sqrt_out = 20'b00010000011101100100;
            11'b00100010000 : sqrt_out = 20'b00010000011111100000;
            11'b00100010001 : sqrt_out = 20'b00010000100001011101;
            11'b00100010010 : sqrt_out = 20'b00010000100011011000;
            11'b00100010011 : sqrt_out = 20'b00010000100101010100;
            11'b00100010100 : sqrt_out = 20'b00010000100111001111;
            11'b00100010101 : sqrt_out = 20'b00010000101001001011;
            11'b00100010110 : sqrt_out = 20'b00010000101011000101;
            11'b00100010111 : sqrt_out = 20'b00010000101101000000;
            11'b00100011000 : sqrt_out = 20'b00010000101110111011;
            11'b00100011001 : sqrt_out = 20'b00010000110000110101;
            11'b00100011010 : sqrt_out = 20'b00010000110010101111;
            11'b00100011011 : sqrt_out = 20'b00010000110100101001;
            11'b00100011100 : sqrt_out = 20'b00010000110110100011;
            11'b00100011101 : sqrt_out = 20'b00010000111000011100;
            11'b00100011110 : sqrt_out = 20'b00010000111010010101;
            11'b00100011111 : sqrt_out = 20'b00010000111100001110;
            11'b00100100000 : sqrt_out = 20'b00010000111110000111;
            11'b00100100001 : sqrt_out = 20'b00010001000000000000;
            11'b00100100010 : sqrt_out = 20'b00010001000001111000;
            11'b00100100011 : sqrt_out = 20'b00010001000011110000;
            11'b00100100100 : sqrt_out = 20'b00010001000101101000;
            11'b00100100101 : sqrt_out = 20'b00010001000111100000;
            11'b00100100110 : sqrt_out = 20'b00010001001001010111;
            11'b00100100111 : sqrt_out = 20'b00010001001011001111;
            11'b00100101000 : sqrt_out = 20'b00010001001101000110;
            11'b00100101001 : sqrt_out = 20'b00010001001110111101;
            11'b00100101010 : sqrt_out = 20'b00010001010000110011;
            11'b00100101011 : sqrt_out = 20'b00010001010010101010;
            11'b00100101100 : sqrt_out = 20'b00010001010100100000;
            11'b00100101101 : sqrt_out = 20'b00010001010110010110;
            11'b00100101110 : sqrt_out = 20'b00010001011000001100;
            11'b00100101111 : sqrt_out = 20'b00010001011010000010;
            11'b00100110000 : sqrt_out = 20'b00010001011011111000;
            11'b00100110001 : sqrt_out = 20'b00010001011101101101;
            11'b00100110010 : sqrt_out = 20'b00010001011111100010;
            11'b00100110011 : sqrt_out = 20'b00010001100001010111;
            11'b00100110100 : sqrt_out = 20'b00010001100011001100;
            11'b00100110101 : sqrt_out = 20'b00010001100101000001;
            11'b00100110110 : sqrt_out = 20'b00010001100110110101;
            11'b00100110111 : sqrt_out = 20'b00010001101000101001;
            11'b00100111000 : sqrt_out = 20'b00010001101010011101;
            11'b00100111001 : sqrt_out = 20'b00010001101100010001;
            11'b00100111010 : sqrt_out = 20'b00010001101110000101;
            11'b00100111011 : sqrt_out = 20'b00010001101111111000;
            11'b00100111100 : sqrt_out = 20'b00010001110001101100;
            11'b00100111101 : sqrt_out = 20'b00010001110011011111;
            11'b00100111110 : sqrt_out = 20'b00010001110101010010;
            11'b00100111111 : sqrt_out = 20'b00010001110111000100;
            11'b00101000000 : sqrt_out = 20'b00010001111000110111;
            11'b00101000001 : sqrt_out = 20'b00010001111010101001;
            11'b00101000010 : sqrt_out = 20'b00010001111100011100;
            11'b00101000011 : sqrt_out = 20'b00010001111110001110;
            11'b00101000100 : sqrt_out = 20'b00010010000000000000;
            11'b00101000101 : sqrt_out = 20'b00010010000001110001;
            11'b00101000110 : sqrt_out = 20'b00010010000011100011;
            11'b00101000111 : sqrt_out = 20'b00010010000101010100;
            11'b00101001000 : sqrt_out = 20'b00010010000111000101;
            11'b00101001001 : sqrt_out = 20'b00010010001000110110;
            11'b00101001010 : sqrt_out = 20'b00010010001010100111;
            11'b00101001011 : sqrt_out = 20'b00010010001100011000;
            11'b00101001100 : sqrt_out = 20'b00010010001110001000;
            11'b00101001101 : sqrt_out = 20'b00010010001111111000;
            11'b00101001110 : sqrt_out = 20'b00010010010001101001;
            11'b00101001111 : sqrt_out = 20'b00010010010011011001;
            11'b00101010000 : sqrt_out = 20'b00010010010101001000;
            11'b00101010001 : sqrt_out = 20'b00010010010110111000;
            11'b00101010010 : sqrt_out = 20'b00010010011000101000;
            11'b00101010011 : sqrt_out = 20'b00010010011010010111;
            11'b00101010100 : sqrt_out = 20'b00010010011100000110;
            11'b00101010101 : sqrt_out = 20'b00010010011101110101;
            11'b00101010110 : sqrt_out = 20'b00010010011111100100;
            11'b00101010111 : sqrt_out = 20'b00010010100001010010;
            11'b00101011000 : sqrt_out = 20'b00010010100011000001;
            11'b00101011001 : sqrt_out = 20'b00010010100100101111;
            11'b00101011010 : sqrt_out = 20'b00010010100110011110;
            11'b00101011011 : sqrt_out = 20'b00010010101000001100;
            11'b00101011100 : sqrt_out = 20'b00010010101001111001;
            11'b00101011101 : sqrt_out = 20'b00010010101011100111;
            11'b00101011110 : sqrt_out = 20'b00010010101101010101;
            11'b00101011111 : sqrt_out = 20'b00010010101111000010;
            11'b00101100000 : sqrt_out = 20'b00010010110000101111;
            11'b00101100001 : sqrt_out = 20'b00010010110010011100;
            11'b00101100010 : sqrt_out = 20'b00010010110100001001;
            11'b00101100011 : sqrt_out = 20'b00010010110101110110;
            11'b00101100100 : sqrt_out = 20'b00010010110111100011;
            11'b00101100101 : sqrt_out = 20'b00010010111001001111;
            11'b00101100110 : sqrt_out = 20'b00010010111010111011;
            11'b00101100111 : sqrt_out = 20'b00010010111100101000;
            11'b00101101000 : sqrt_out = 20'b00010010111110010100;
            11'b00101101001 : sqrt_out = 20'b00010011000000000000;
            11'b00101101010 : sqrt_out = 20'b00010011000001101011;
            11'b00101101011 : sqrt_out = 20'b00010011000011010111;
            11'b00101101100 : sqrt_out = 20'b00010011000101000010;
            11'b00101101101 : sqrt_out = 20'b00010011000110101101;
            11'b00101101110 : sqrt_out = 20'b00010011001000011001;
            11'b00101101111 : sqrt_out = 20'b00010011001010000100;
            11'b00101110000 : sqrt_out = 20'b00010011001011101110;
            11'b00101110001 : sqrt_out = 20'b00010011001101011001;
            11'b00101110010 : sqrt_out = 20'b00010011001111000100;
            11'b00101110011 : sqrt_out = 20'b00010011010000101110;
            11'b00101110100 : sqrt_out = 20'b00010011010010011000;
            11'b00101110101 : sqrt_out = 20'b00010011010100000010;
            11'b00101110110 : sqrt_out = 20'b00010011010101101100;
            11'b00101110111 : sqrt_out = 20'b00010011010111010110;
            11'b00101111000 : sqrt_out = 20'b00010011011001000000;
            11'b00101111001 : sqrt_out = 20'b00010011011010101001;
            11'b00101111010 : sqrt_out = 20'b00010011011100010011;
            11'b00101111011 : sqrt_out = 20'b00010011011101111100;
            11'b00101111100 : sqrt_out = 20'b00010011011111100101;
            11'b00101111101 : sqrt_out = 20'b00010011100001001110;
            11'b00101111110 : sqrt_out = 20'b00010011100010110111;
            11'b00101111111 : sqrt_out = 20'b00010011100100100000;
            11'b00110000000 : sqrt_out = 20'b00010011100110001000;
            11'b00110000001 : sqrt_out = 20'b00010011100111110001;
            11'b00110000010 : sqrt_out = 20'b00010011101001011001;
            11'b00110000011 : sqrt_out = 20'b00010011101011000001;
            11'b00110000100 : sqrt_out = 20'b00010011101100101001;
            11'b00110000101 : sqrt_out = 20'b00010011101110010001;
            11'b00110000110 : sqrt_out = 20'b00010011101111111001;
            11'b00110000111 : sqrt_out = 20'b00010011110001100001;
            11'b00110001000 : sqrt_out = 20'b00010011110011001000;
            11'b00110001001 : sqrt_out = 20'b00010011110100110000;
            11'b00110001010 : sqrt_out = 20'b00010011110110010111;
            11'b00110001011 : sqrt_out = 20'b00010011110111111110;
            11'b00110001100 : sqrt_out = 20'b00010011111001100101;
            11'b00110001101 : sqrt_out = 20'b00010011111011001100;
            11'b00110001110 : sqrt_out = 20'b00010011111100110010;
            11'b00110001111 : sqrt_out = 20'b00010011111110011001;
            11'b00110010000 : sqrt_out = 20'b00010100000000000000;
            11'b00110010001 : sqrt_out = 20'b00010100000001100110;
            11'b00110010010 : sqrt_out = 20'b00010100000011001100;
            11'b00110010011 : sqrt_out = 20'b00010100000100110010;
            11'b00110010100 : sqrt_out = 20'b00010100000110011000;
            11'b00110010101 : sqrt_out = 20'b00010100000111111110;
            11'b00110010110 : sqrt_out = 20'b00010100001001100100;
            11'b00110010111 : sqrt_out = 20'b00010100001011001001;
            11'b00110011000 : sqrt_out = 20'b00010100001100101111;
            11'b00110011001 : sqrt_out = 20'b00010100001110010100;
            11'b00110011010 : sqrt_out = 20'b00010100001111111001;
            11'b00110011011 : sqrt_out = 20'b00010100010001011110;
            11'b00110011100 : sqrt_out = 20'b00010100010011000011;
            11'b00110011101 : sqrt_out = 20'b00010100010100101000;
            11'b00110011110 : sqrt_out = 20'b00010100010110001101;
            11'b00110011111 : sqrt_out = 20'b00010100010111110001;
            11'b00110100000 : sqrt_out = 20'b00010100011001010110;
            11'b00110100001 : sqrt_out = 20'b00010100011010111010;
            11'b00110100010 : sqrt_out = 20'b00010100011100011110;
            11'b00110100011 : sqrt_out = 20'b00010100011110000011;
            11'b00110100100 : sqrt_out = 20'b00010100011111100111;
            11'b00110100101 : sqrt_out = 20'b00010100100001001010;
            11'b00110100110 : sqrt_out = 20'b00010100100010101110;
            11'b00110100111 : sqrt_out = 20'b00010100100100010010;
            11'b00110101000 : sqrt_out = 20'b00010100100101110101;
            11'b00110101001 : sqrt_out = 20'b00010100100111011001;
            11'b00110101010 : sqrt_out = 20'b00010100101000111100;
            11'b00110101011 : sqrt_out = 20'b00010100101010011111;
            11'b00110101100 : sqrt_out = 20'b00010100101100000010;
            11'b00110101101 : sqrt_out = 20'b00010100101101100101;
            11'b00110101110 : sqrt_out = 20'b00010100101111001000;
            11'b00110101111 : sqrt_out = 20'b00010100110000101011;
            11'b00110110000 : sqrt_out = 20'b00010100110010001101;
            11'b00110110001 : sqrt_out = 20'b00010100110011110000;
            11'b00110110010 : sqrt_out = 20'b00010100110101010010;
            11'b00110110011 : sqrt_out = 20'b00010100110110110100;
            11'b00110110100 : sqrt_out = 20'b00010100111000010110;
            11'b00110110101 : sqrt_out = 20'b00010100111001111001;
            11'b00110110110 : sqrt_out = 20'b00010100111011011010;
            11'b00110110111 : sqrt_out = 20'b00010100111100111100;
            11'b00110111000 : sqrt_out = 20'b00010100111110011110;
            11'b00110111001 : sqrt_out = 20'b00010101000000000000;
            11'b00110111010 : sqrt_out = 20'b00010101000001100001;
            11'b00110111011 : sqrt_out = 20'b00010101000011000010;
            11'b00110111100 : sqrt_out = 20'b00010101000100100100;
            11'b00110111101 : sqrt_out = 20'b00010101000110000101;
            11'b00110111110 : sqrt_out = 20'b00010101000111100110;
            11'b00110111111 : sqrt_out = 20'b00010101001001000111;
            11'b00111000000 : sqrt_out = 20'b00010101001010100111;
            11'b00111000001 : sqrt_out = 20'b00010101001100001000;
            11'b00111000010 : sqrt_out = 20'b00010101001101101001;
            11'b00111000011 : sqrt_out = 20'b00010101001111001001;
            11'b00111000100 : sqrt_out = 20'b00010101010000101010;
            11'b00111000101 : sqrt_out = 20'b00010101010010001010;
            11'b00111000110 : sqrt_out = 20'b00010101010011101010;
            11'b00111000111 : sqrt_out = 20'b00010101010101001010;
            11'b00111001000 : sqrt_out = 20'b00010101010110101010;
            11'b00111001001 : sqrt_out = 20'b00010101011000001010;
            11'b00111001010 : sqrt_out = 20'b00010101011001101010;
            11'b00111001011 : sqrt_out = 20'b00010101011011001001;
            11'b00111001100 : sqrt_out = 20'b00010101011100101001;
            11'b00111001101 : sqrt_out = 20'b00010101011110001000;
            11'b00111001110 : sqrt_out = 20'b00010101011111101000;
            11'b00111001111 : sqrt_out = 20'b00010101100001000111;
            11'b00111010000 : sqrt_out = 20'b00010101100010100110;
            11'b00111010001 : sqrt_out = 20'b00010101100100000101;
            11'b00111010010 : sqrt_out = 20'b00010101100101100100;
            11'b00111010011 : sqrt_out = 20'b00010101100111000011;
            11'b00111010100 : sqrt_out = 20'b00010101101000100010;
            11'b00111010101 : sqrt_out = 20'b00010101101010000000;
            11'b00111010110 : sqrt_out = 20'b00010101101011011111;
            11'b00111010111 : sqrt_out = 20'b00010101101100111101;
            11'b00111011000 : sqrt_out = 20'b00010101101110011011;
            11'b00111011001 : sqrt_out = 20'b00010101101111111010;
            11'b00111011010 : sqrt_out = 20'b00010101110001011000;
            11'b00111011011 : sqrt_out = 20'b00010101110010110110;
            11'b00111011100 : sqrt_out = 20'b00010101110100010100;
            11'b00111011101 : sqrt_out = 20'b00010101110101110001;
            11'b00111011110 : sqrt_out = 20'b00010101110111001111;
            11'b00111011111 : sqrt_out = 20'b00010101111000101101;
            11'b00111100000 : sqrt_out = 20'b00010101111010001010;
            11'b00111100001 : sqrt_out = 20'b00010101111011101000;
            11'b00111100010 : sqrt_out = 20'b00010101111101000101;
            11'b00111100011 : sqrt_out = 20'b00010101111110100010;
            11'b00111100100 : sqrt_out = 20'b00010110000000000000;
            11'b00111100101 : sqrt_out = 20'b00010110000001011101;
            11'b00111100110 : sqrt_out = 20'b00010110000010111001;
            11'b00111100111 : sqrt_out = 20'b00010110000100010110;
            11'b00111101000 : sqrt_out = 20'b00010110000101110011;
            11'b00111101001 : sqrt_out = 20'b00010110000111010000;
            11'b00111101010 : sqrt_out = 20'b00010110001000101100;
            11'b00111101011 : sqrt_out = 20'b00010110001010001001;
            11'b00111101100 : sqrt_out = 20'b00010110001011100101;
            11'b00111101101 : sqrt_out = 20'b00010110001101000001;
            11'b00111101110 : sqrt_out = 20'b00010110001110011110;
            11'b00111101111 : sqrt_out = 20'b00010110001111111010;
            11'b00111110000 : sqrt_out = 20'b00010110010001010110;
            11'b00111110001 : sqrt_out = 20'b00010110010010110010;
            11'b00111110010 : sqrt_out = 20'b00010110010100001101;
            11'b00111110011 : sqrt_out = 20'b00010110010101101001;
            11'b00111110100 : sqrt_out = 20'b00010110010111000101;
            11'b00111110101 : sqrt_out = 20'b00010110011000100000;
            11'b00111110110 : sqrt_out = 20'b00010110011001111100;
            11'b00111110111 : sqrt_out = 20'b00010110011011010111;
            11'b00111111000 : sqrt_out = 20'b00010110011100110010;
            11'b00111111001 : sqrt_out = 20'b00010110011110001110;
            11'b00111111010 : sqrt_out = 20'b00010110011111101001;
            11'b00111111011 : sqrt_out = 20'b00010110100001000100;
            11'b00111111100 : sqrt_out = 20'b00010110100010011111;
            11'b00111111101 : sqrt_out = 20'b00010110100011111001;
            11'b00111111110 : sqrt_out = 20'b00010110100101010100;
            11'b00111111111 : sqrt_out = 20'b00010110100110101111;


            11'b00010000000 : sqrt_out = 20'b00001011010100000100;
            11'b00010000001 : sqrt_out = 20'b00001011010110111001;
            11'b00010000010 : sqrt_out = 20'b00001011011001101101;
            11'b00010000011 : sqrt_out = 20'b00001011011100100000;
            11'b00010000100 : sqrt_out = 20'b00001011011111010011;
            11'b00010000101 : sqrt_out = 20'b00001011100010000101;
            11'b00010000110 : sqrt_out = 20'b00001011100100110110;
            11'b00010000111 : sqrt_out = 20'b00001011100111100111;
            11'b00010001000 : sqrt_out = 20'b00001011101010010111;
            11'b00010001001 : sqrt_out = 20'b00001011101101000110;
            11'b00010001010 : sqrt_out = 20'b00001011101111110101;
            11'b00010001011 : sqrt_out = 20'b00001011110010100011;
            11'b00010001100 : sqrt_out = 20'b00001011110101010000;
            11'b00010001101 : sqrt_out = 20'b00001011110111111101;
            11'b00010001110 : sqrt_out = 20'b00001011111010101001;
            11'b00010001111 : sqrt_out = 20'b00001011111101010101;
            11'b00010010000 : sqrt_out = 20'b00001100000000000000;
            11'b00010010001 : sqrt_out = 20'b00001100000010101010;
            11'b00010010010 : sqrt_out = 20'b00001100000101010100;
            11'b00010010011 : sqrt_out = 20'b00001100000111111101;
            11'b00010010100 : sqrt_out = 20'b00001100001010100101;
            11'b00010010101 : sqrt_out = 20'b00001100001101001110;
            11'b00010010110 : sqrt_out = 20'b00001100001111110101;
            11'b00010010111 : sqrt_out = 20'b00001100010010011100;
            11'b00010011000 : sqrt_out = 20'b00001100010101000010;
            11'b00010011001 : sqrt_out = 20'b00001100010111101000;
            11'b00010011010 : sqrt_out = 20'b00001100011010001110;
            11'b00010011011 : sqrt_out = 20'b00001100011100110010;
            11'b00010011100 : sqrt_out = 20'b00001100011111010111;
            11'b00010011101 : sqrt_out = 20'b00001100100001111010;
            11'b00010011110 : sqrt_out = 20'b00001100100100011101;
            11'b00010011111 : sqrt_out = 20'b00001100100111000000;
            11'b00010100000 : sqrt_out = 20'b00001100101001100010;
            11'b00010100001 : sqrt_out = 20'b00001100101100000100;
            11'b00010100010 : sqrt_out = 20'b00001100101110100101;
            11'b00010100011 : sqrt_out = 20'b00001100110001000110;
            11'b00010100100 : sqrt_out = 20'b00001100110011100110;
            11'b00010100101 : sqrt_out = 20'b00001100110110000110;
            11'b00010100110 : sqrt_out = 20'b00001100111000100101;
            11'b00010100111 : sqrt_out = 20'b00001100111011000011;
            11'b00010101000 : sqrt_out = 20'b00001100111101100010;
            11'b00010101001 : sqrt_out = 20'b00001101000000000000;
            11'b00010101010 : sqrt_out = 20'b00001101000010011101;
            11'b00010101011 : sqrt_out = 20'b00001101000100111010;
            11'b00010101100 : sqrt_out = 20'b00001101000111010110;
            11'b00010101101 : sqrt_out = 20'b00001101001001110010;
            11'b00010101110 : sqrt_out = 20'b00001101001100001101;
            11'b00010101111 : sqrt_out = 20'b00001101001110101000;
            11'b00010110000 : sqrt_out = 20'b00001101010001000011;
            11'b00010110001 : sqrt_out = 20'b00001101010011011101;
            11'b00010110010 : sqrt_out = 20'b00001101010101110111;
            11'b00010110011 : sqrt_out = 20'b00001101011000010000;
            11'b00010110100 : sqrt_out = 20'b00001101011010101001;
            11'b00010110101 : sqrt_out = 20'b00001101011101000010;
            11'b00010110110 : sqrt_out = 20'b00001101011111011010;
            11'b00010110111 : sqrt_out = 20'b00001101100001110001;
            11'b00010111000 : sqrt_out = 20'b00001101100100001000;
            11'b00010111001 : sqrt_out = 20'b00001101100110011111;
            11'b00010111010 : sqrt_out = 20'b00001101101000110101;
            11'b00010111011 : sqrt_out = 20'b00001101101011001011;
            11'b00010111100 : sqrt_out = 20'b00001101101101100001;
            11'b00010111101 : sqrt_out = 20'b00001101101111110110;
            11'b00010111110 : sqrt_out = 20'b00001101110010001011;
            11'b00010111111 : sqrt_out = 20'b00001101110100011111;
            11'b00011000000 : sqrt_out = 20'b00001101110110110011;
            11'b00011000001 : sqrt_out = 20'b00001101111001000111;
            11'b00011000010 : sqrt_out = 20'b00001101111011011010;
            11'b00011000011 : sqrt_out = 20'b00001101111101101101;
            11'b00011000100 : sqrt_out = 20'b00001110000000000000;
            11'b00011000101 : sqrt_out = 20'b00001110000010010010;
            11'b00011000110 : sqrt_out = 20'b00001110000100100011;
            11'b00011000111 : sqrt_out = 20'b00001110000110110101;
            11'b00011001000 : sqrt_out = 20'b00001110001001000110;
            11'b00011001001 : sqrt_out = 20'b00001110001011010110;
            11'b00011001010 : sqrt_out = 20'b00001110001101100111;
            11'b00011001011 : sqrt_out = 20'b00001110001111110111;
            11'b00011001100 : sqrt_out = 20'b00001110010010000110;
            11'b00011001101 : sqrt_out = 20'b00001110010100010101;
            11'b00011001110 : sqrt_out = 20'b00001110010110100100;
            11'b00011001111 : sqrt_out = 20'b00001110011000110011;
            11'b00011010000 : sqrt_out = 20'b00001110011011000001;
            11'b00011010001 : sqrt_out = 20'b00001110011101001111;
            11'b00011010010 : sqrt_out = 20'b00001110011111011100;
            11'b00011010011 : sqrt_out = 20'b00001110100001101001;
            11'b00011010100 : sqrt_out = 20'b00001110100011110110;
            11'b00011010101 : sqrt_out = 20'b00001110100110000011;
            11'b00011010110 : sqrt_out = 20'b00001110101000001111;
            11'b00011010111 : sqrt_out = 20'b00001110101010011011;
            11'b00011011000 : sqrt_out = 20'b00001110101100100110;
            11'b00011011001 : sqrt_out = 20'b00001110101110110001;
            11'b00011011010 : sqrt_out = 20'b00001110110000111100;
            11'b00011011011 : sqrt_out = 20'b00001110110011000111;
            11'b00011011100 : sqrt_out = 20'b00001110110101010001;
            11'b00011011101 : sqrt_out = 20'b00001110110111011011;
            11'b00011011110 : sqrt_out = 20'b00001110111001100101;
            11'b00011011111 : sqrt_out = 20'b00001110111011101110;
            11'b00011100000 : sqrt_out = 20'b00001110111101110111;
            11'b00011100001 : sqrt_out = 20'b00001111000000000000;
            11'b00011100010 : sqrt_out = 20'b00001111000010001000;
            11'b00011100011 : sqrt_out = 20'b00001111000100010000;
            11'b00011100100 : sqrt_out = 20'b00001111000110011000;
            11'b00011100101 : sqrt_out = 20'b00001111001000011111;
            11'b00011100110 : sqrt_out = 20'b00001111001010100110;
            11'b00011100111 : sqrt_out = 20'b00001111001100101101;
            11'b00011101000 : sqrt_out = 20'b00001111001110110100;
            11'b00011101001 : sqrt_out = 20'b00001111010000111010;
            11'b00011101010 : sqrt_out = 20'b00001111010011000000;
            11'b00011101011 : sqrt_out = 20'b00001111010101000110;
            11'b00011101100 : sqrt_out = 20'b00001111010111001011;
            11'b00011101101 : sqrt_out = 20'b00001111011001010001;
            11'b00011101110 : sqrt_out = 20'b00001111011011010110;
            11'b00011101111 : sqrt_out = 20'b00001111011101011010;
            11'b00011110000 : sqrt_out = 20'b00001111011111011110;
            11'b00011110001 : sqrt_out = 20'b00001111100001100011;
            11'b00011110010 : sqrt_out = 20'b00001111100011100110;
            11'b00011110011 : sqrt_out = 20'b00001111100101101010;
            11'b00011110100 : sqrt_out = 20'b00001111100111101101;
            11'b00011110101 : sqrt_out = 20'b00001111101001110000;
            11'b00011110110 : sqrt_out = 20'b00001111101011110011;
            11'b00011110111 : sqrt_out = 20'b00001111101101110101;
            11'b00011111000 : sqrt_out = 20'b00001111101111110111;
            11'b00011111001 : sqrt_out = 20'b00001111110001111001;
            11'b00011111010 : sqrt_out = 20'b00001111110011111011;
            11'b00011111011 : sqrt_out = 20'b00001111110101111100;
            11'b00011111100 : sqrt_out = 20'b00001111110111111101;
            11'b00011111101 : sqrt_out = 20'b00001111111001111110;
            11'b00011111110 : sqrt_out = 20'b00001111111011111111;
            11'b00011111111 : sqrt_out = 20'b00001111111101111111;
            
            11'b00001000000 : sqrt_out = 20'b00001000000000000000;
            11'b00001000001 : sqrt_out = 20'b00001000000011111111;
            11'b00001000010 : sqrt_out = 20'b00001000000111111100;
            11'b00001000011 : sqrt_out = 20'b00001000001011110111;
            11'b00001000100 : sqrt_out = 20'b00001000001111110000;
            11'b00001000101 : sqrt_out = 20'b00001000010011100111;
            11'b00001000110 : sqrt_out = 20'b00001000010111011101;
            11'b00001000111 : sqrt_out = 20'b00001000011011010001;
            11'b00001001000 : sqrt_out = 20'b00001000011111000011;
            11'b00001001001 : sqrt_out = 20'b00001000100010110100;
            11'b00001001010 : sqrt_out = 20'b00001000100110100011;
            11'b00001001011 : sqrt_out = 20'b00001000101010010000;
            11'b00001001100 : sqrt_out = 20'b00001000101101111100;
            11'b00001001101 : sqrt_out = 20'b00001000110001100110;
            11'b00001001110 : sqrt_out = 20'b00001000110101001110;
            11'b00001001111 : sqrt_out = 20'b00001000111000110110;
            11'b00001010000 : sqrt_out = 20'b00001000111100011011;
            11'b00001010001 : sqrt_out = 20'b00001001000000000000;
            11'b00001010010 : sqrt_out = 20'b00001001000011100010;
            11'b00001010011 : sqrt_out = 20'b00001001000111000100;
            11'b00001010100 : sqrt_out = 20'b00001001001010100100;
            11'b00001010101 : sqrt_out = 20'b00001001001110000011;
            11'b00001010110 : sqrt_out = 20'b00001001010001100000;
            11'b00001010111 : sqrt_out = 20'b00001001010100111100;
            11'b00001011000 : sqrt_out = 20'b00001001011000010111;
            11'b00001011001 : sqrt_out = 20'b00001001011011110001;
            11'b00001011010 : sqrt_out = 20'b00001001011111001010;
            11'b00001011011 : sqrt_out = 20'b00001001100010100001;
            11'b00001011100 : sqrt_out = 20'b00001001100101110111;
            11'b00001011101 : sqrt_out = 20'b00001001101001001100;
            11'b00001011110 : sqrt_out = 20'b00001001101100100000;
            11'b00001011111 : sqrt_out = 20'b00001001101111110010;
            11'b00001100000 : sqrt_out = 20'b00001001110011000100;
            11'b00001100001 : sqrt_out = 20'b00001001110110010100;
            11'b00001100010 : sqrt_out = 20'b00001001111001100100;
            11'b00001100011 : sqrt_out = 20'b00001001111100110010;
            11'b00001100100 : sqrt_out = 20'b00001010000000000000;
            11'b00001100101 : sqrt_out = 20'b00001010000011001100;
            11'b00001100110 : sqrt_out = 20'b00001010000110010111;
            11'b00001100111 : sqrt_out = 20'b00001010001001100001;
            11'b00001101000 : sqrt_out = 20'b00001010001100101011;
            11'b00001101001 : sqrt_out = 20'b00001010001111110011;
            11'b00001101010 : sqrt_out = 20'b00001010010010111010;
            11'b00001101011 : sqrt_out = 20'b00001010010110000001;
            11'b00001101100 : sqrt_out = 20'b00001010011001000110;
            11'b00001101101 : sqrt_out = 20'b00001010011100001011;
            11'b00001101110 : sqrt_out = 20'b00001010011111001111;
            11'b00001101111 : sqrt_out = 20'b00001010100010010010;
            11'b00001110000 : sqrt_out = 20'b00001010100101010011;
            11'b00001110001 : sqrt_out = 20'b00001010101000010101;
            11'b00001110010 : sqrt_out = 20'b00001010101011010101;
            11'b00001110011 : sqrt_out = 20'b00001010101110010100;
            11'b00001110100 : sqrt_out = 20'b00001010110001010011;
            11'b00001110101 : sqrt_out = 20'b00001010110100010001;
            11'b00001110110 : sqrt_out = 20'b00001010110111001101;
            11'b00001110111 : sqrt_out = 20'b00001010111010001010;
            11'b00001111000 : sqrt_out = 20'b00001010111101000101;
            11'b00001111001 : sqrt_out = 20'b00001011000000000000;
            11'b00001111010 : sqrt_out = 20'b00001011000010111001;
            11'b00001111011 : sqrt_out = 20'b00001011000101110010;
            11'b00001111100 : sqrt_out = 20'b00001011001000101011;
            11'b00001111101 : sqrt_out = 20'b00001011001011100010;
            11'b00001111110 : sqrt_out = 20'b00001011001110011001;
            11'b00001111111 : sqrt_out = 20'b00001011010001001111;

            11'b00000100000 : sqrt_out = 20'b00000101101010000010;
            11'b00000100001 : sqrt_out = 20'b00000101101111101001;
            11'b00000100010 : sqrt_out = 20'b00000101110101001011;
            11'b00000100011 : sqrt_out = 20'b00000101111010101000;
            11'b00000100100 : sqrt_out = 20'b00000110000000000000;
            11'b00000100101 : sqrt_out = 20'b00000110000101010010;
            11'b00000100110 : sqrt_out = 20'b00000110001010100001;
            11'b00000100111 : sqrt_out = 20'b00000110001111101011;
            11'b00000101000 : sqrt_out = 20'b00000110010100110001;
            11'b00000101001 : sqrt_out = 20'b00000110011001110011;
            11'b00000101010 : sqrt_out = 20'b00000110011110110001;
            11'b00000101011 : sqrt_out = 20'b00000110100011101011;
            11'b00000101100 : sqrt_out = 20'b00000110101000100001;
            11'b00000101101 : sqrt_out = 20'b00000110101101010100;
            11'b00000101110 : sqrt_out = 20'b00000110110010000100;
            11'b00000101111 : sqrt_out = 20'b00000110110110110000;
            11'b00000110000 : sqrt_out = 20'b00000110111011011001;
            11'b00000110001 : sqrt_out = 20'b00000111000000000000;
            11'b00000110010 : sqrt_out = 20'b00000111000100100011;
            11'b00000110011 : sqrt_out = 20'b00000111001001000011;
            11'b00000110100 : sqrt_out = 20'b00000111001101100000;
            11'b00000110101 : sqrt_out = 20'b00000111010001111011;
            11'b00000110110 : sqrt_out = 20'b00000111010110010011;
            11'b00000110111 : sqrt_out = 20'b00000111011010101000;
            11'b00000111000 : sqrt_out = 20'b00000111011110111011;
            11'b00000111001 : sqrt_out = 20'b00000111100011001100;
            11'b00000111010 : sqrt_out = 20'b00000111100111011010;
            11'b00000111011 : sqrt_out = 20'b00000111101011100101;
            11'b00000111100 : sqrt_out = 20'b00000111101111101111;
            11'b00000111101 : sqrt_out = 20'b00000111110011110110;
            11'b00000111110 : sqrt_out = 20'b00000111110111111011;
            11'b00000111111 : sqrt_out = 20'b00000111111011111110;

            11'b00000010000 : sqrt_out = 20'b00000100000000000000;
            11'b00000010001 : sqrt_out = 20'b00000100000111111000;
            11'b00000010010 : sqrt_out = 20'b00000100001111100001;
            11'b00000010011 : sqrt_out = 20'b00000100010110111110;
            11'b00000010100 : sqrt_out = 20'b00000100011110001101;
            11'b00000010101 : sqrt_out = 20'b00000100100101010010;
            11'b00000010110 : sqrt_out = 20'b00000100101100001011;
            11'b00000010111 : sqrt_out = 20'b00000100110010111011;
            11'b00000011000 : sqrt_out = 20'b00000100111001100010;
            11'b00000011001 : sqrt_out = 20'b00000101000000000000;
            11'b00000011010 : sqrt_out = 20'b00000101000110010101;
            11'b00000011011 : sqrt_out = 20'b00000101001100100011;
            11'b00000011100 : sqrt_out = 20'b00000101010010101001;
            11'b00000011101 : sqrt_out = 20'b00000101011000101001;
            11'b00000011110 : sqrt_out = 20'b00000101011110100010;
            11'b00000011111 : sqrt_out = 20'b00000101100100010101;
            11'b00000001000 : sqrt_out = 20'b00000010110101000001;
            11'b00000001001 : sqrt_out = 20'b00000011000000000000;
            11'b00000001010 : sqrt_out = 20'b00000011001010011000;
            11'b00000001011 : sqrt_out = 20'b00000011010100010000;
            11'b00000001100 : sqrt_out = 20'b00000011011101101100;
            11'b00000001101 : sqrt_out = 20'b00000011100110110000;
            11'b00000001110 : sqrt_out = 20'b00000011101111011101;
            11'b00000001111 : sqrt_out = 20'b00000011110111110111;
            11'b00000000100 : sqrt_out = 20'b00000010000000000000;
            11'b00000000101 : sqrt_out = 20'b00000010001111000110;
            11'b00000000110 : sqrt_out = 20'b00000010011100110001;
            11'b00000000111 : sqrt_out = 20'b00000010101001010100;
            11'b00000000010 : sqrt_out = 20'b00000001011010100000;
            11'b00000000011 : sqrt_out = 20'b00000001101110110110;

            11'b00000000001 : sqrt_out = 20'b00000001000000000000;

        endcase
    end
endmodule